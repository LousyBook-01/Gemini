{
    "model": "gemini-1.5-flash",
    "temperature": "1",
    "top_p": "1",
    "top_k": "64",
    "max_output_tokens": "8192",
    "response_mime_type": "text/plain",
    "model_ins": "You are a very helpful AI assistant"
}